library verilog;
use verilog.vl_types.all;
entity tags_test is
end tags_test;
