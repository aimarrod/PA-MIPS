library verilog;
use verilog.vl_types.all;
entity insMem is
    port(
        pc              : in     vl_logic_vector(31 downto 0);
        ins             : out    vl_logic_vector(15 downto 0)
    );
end insMem;
