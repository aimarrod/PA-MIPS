library verilog;
use verilog.vl_types.all;
entity reorder_buffer is
    port(
        clk             : in     vl_logic;
        stall           : in     vl_logic;
        alu             : in     vl_logic_vector(2 downto 0);
        alu_we          : in     vl_logic;
        alu_rd          : in     vl_logic_vector(4 downto 0);
        alu_pc          : in     vl_logic_vector(31 downto 0);
        alu_ex          : in     vl_logic;
        alu_val         : in     vl_logic_vector(31 downto 0);
        alu_store       : in     vl_logic;
        alu_addr        : in     vl_logic_vector(31 downto 0);
        alu_pass        : in     vl_logic;
        load            : in     vl_logic_vector(2 downto 0);
        load_pc         : in     vl_logic_vector(31 downto 0);
        load_we         : in     vl_logic;
        load_rd         : in     vl_logic_vector(4 downto 0);
        load_ex         : in     vl_logic;
        load_val        : in     vl_logic_vector(31 downto 0);
        load_addr       : in     vl_logic_vector(31 downto 0);
        slow            : in     vl_logic_vector(2 downto 0);
        slow_we         : in     vl_logic;
        slow_pc         : in     vl_logic_vector(31 downto 0);
        slow_rd         : in     vl_logic_vector(4 downto 0);
        slow_ex         : in     vl_logic;
        slow_val        : in     vl_logic_vector(31 downto 0);
        val_out         : out    vl_logic_vector(31 downto 0);
        rd_out          : out    vl_logic_vector(4 downto 0);
        we              : out    vl_logic;
        ex_out          : out    vl_logic;
        store_out       : out    vl_logic;
        pc_out          : out    vl_logic_vector(31 downto 0);
        addr_out        : out    vl_logic_vector(31 downto 0);
        stores          : out    vl_logic;
        tail_out        : out    vl_logic_vector(2 downto 0);
        next_head       : in     vl_logic;
        destination_0   : out    vl_logic_vector(4 downto 0);
        destination_1   : out    vl_logic_vector(4 downto 0);
        destination_2   : out    vl_logic_vector(4 downto 0);
        destination_3   : out    vl_logic_vector(4 downto 0);
        destination_4   : out    vl_logic_vector(4 downto 0);
        destination_5   : out    vl_logic_vector(4 downto 0);
        destination_6   : out    vl_logic_vector(4 downto 0);
        destination_7   : out    vl_logic_vector(4 downto 0);
        val_0           : out    vl_logic_vector(31 downto 0);
        val_1           : out    vl_logic_vector(31 downto 0);
        val_2           : out    vl_logic_vector(31 downto 0);
        val_3           : out    vl_logic_vector(31 downto 0);
        val_4           : out    vl_logic_vector(31 downto 0);
        val_5           : out    vl_logic_vector(31 downto 0);
        val_6           : out    vl_logic_vector(31 downto 0);
        val_7           : out    vl_logic_vector(31 downto 0);
        valids          : out    vl_logic_vector(7 downto 0)
    );
end reorder_buffer;
